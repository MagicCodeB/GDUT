//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Dec 26 13:11:21 2020
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// Zhq
module Zhq(
    // Inputs
    DataIn,
    // Outputs
    bai,
    ge,
    shi
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [7:0] DataIn;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [3:0] bai;
output [3:0] ge;
output [3:0] shi;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [3:0] bai_net_0;
wire   [7:0] DataIn;
wire   [3:0] ge_net_0;
wire   [3:0] shi_net_0;
wire   [3:0] ge_net_1;
wire   [3:0] shi_net_1;
wire   [3:0] bai_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign ge_net_1  = ge_net_0;
assign ge[3:0]   = ge_net_1;
assign shi_net_1 = shi_net_0;
assign shi[3:0]  = shi_net_1;
assign bai_net_1 = bai_net_0;
assign bai[3:0]  = bai_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------W_zh5
W_zh5 W_zh5_0(
        // Inputs
        .DataIn ( DataIn ),
        // Outputs
        .ge     ( ge_net_0 ),
        .shi    ( shi_net_0 ),
        .bai    ( bai_net_0 ) 
        );


endmodule
